module char_rom #(
    parameter DATA_WIDTH = 35,     // Width of ROM data (35 bits for each character)
    parameter ADDR_WIDTH = 7,      // Address width
    parameter ADDR_MIN = 32,
    parameter ADDR_MAX = 127
)(
    input wire [ADDR_WIDTH-1:0] address,
    output wire [DATA_WIDTH-1:0] data
);

reg [DATA_WIDTH-1:0] d;

assign data = { d[2], d[24], d[11], d[23], d[33], d[34], d[30], d[9], d[4], d[16], d[22], d[17], d[20], d[8], d[29], d[3], d[25], d[10], d[32], d[1], d[19], d[14], d[7], d[13], d[28], d[21], d[15], d[5], d[6], d[0], d[31], d[18], d[27], d[12], d[26] };

reg [DATA_WIDTH-1:0] mem [0:ADDR_MAX-ADDR_MIN];

initial begin
    $readmemb("font.bin", mem);  // load char bitmaps from file
end

assign d = |address[ADDR_WIDTH-1:5] ? mem[address-ADDR_MIN] : '1;

endmodule
